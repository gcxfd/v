#!/usr/bin/env v run

module main

fn main() {
	println('Hello World!')
}
