#!/usr/bin/env -S v run

module main

fn main() {
	println('Hello World!')
}
